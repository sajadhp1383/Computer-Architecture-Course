module Rat_Controller(input clk, rst, start, run, cout, invalid, finish, empty1, empty2, full1, full2,
                        output logic ldC, ldX, ldY, Izc, SelMux5, DinMem, push1, pop1, push2, pop2,
                            cen, WR, RD, fail, done);


endmodule