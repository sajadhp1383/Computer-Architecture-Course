module datapath();

    

endmodule