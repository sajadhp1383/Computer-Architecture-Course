library verilog;
use verilog.vl_types.all;
entity TEST_RISCV is
end TEST_RISCV;
